----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 22.12.2020 19:05:42
-- Design Name: 
-- Module Name: memory - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity memory is
  Port ( address: in std_logic_vector (31 downto 0);
        write_data: in std_logic_vector (31 downto 0);
        clk: in std_logic;
        MW: in std_logic;
        read_data: out std_logic_vector (31 downto 0) );
end memory;

architecture Behavioral of memory is

    -- we will use the least significant 9 bit of the address – array(0 to 512)
    type mem_array is array(0 to 511) of std_logic_vector(31 downto 0);

    begin mem_process: process (address, write_data, clk, MW)
    
    variable data_mem: mem_array :=(
    
       -- ZEROETH SET
       
       
       -- start and load all the registers with different values
       X"00000000",
       
       -- opcode = 00000000000000000, dr = 00000, sa = 00000,  sb = 00011
       -- reg 0
       X"00000003",
       
       -- opcode = 00000000000000000, dr = 00001, sa = 00000,  sb = 00011
       -- reg 1
       X"00000402",
       
       -- opcode = 00000000000000000, dr = 00010, sa = 00000,  sb = 00001
       -- reg 2
       X"00000801",
       
       -- opcode = 00000000000000000, dr = 00011, sa = 00000,  sb = 00000
       -- reg 3
       X"00000C00",
       
       -- opcode = 00000000000000000, dr = 00100, sa = 00000,  sb = 00011
       -- reg 4
       X"00001003",
       
       -- opcode = 00000000000000000, dr = 00101, sa = 00000,  sb = 00010
       -- reg 5
       X"00001402",
       
       -- opcode = 00000000000000000, dr = 00110, sa = 00000,  sb = 00001
       -- reg 6
       X"00001801",
       
       -- opcode = 00000000000000000, dr = 00111, sa = 00000,  sb = 00000
       -- reg 7
       X"00001C00",
       
       -- opcode = 00000000000000000, dr = 01000, sa = 00000,  sb = 00011
       -- reg 8
       X"00002003",
       
       -- opcode = 00000000000000000, dr = 01001, sa = 00000,  sb = 00011
       -- reg 9
       X"00002402",
       
       -- opcode = 00000000000000000, dr = 01010, sa = 00000,  sb = 00001
       -- reg 10
       X"00002801",
       
       -- opcode = 00000000000000000, dr = 01011, sa = 00000,  sb = 00000
       -- reg 11
       X"00002C00",
       
       -- opcode = 00000000000000000, dr = 01100, sa = 00000,  sb = 00011
       -- reg 12
       X"00003003",
       
       -- opcode = 00000000000000000, dr = 01101, sa = 00000,  sb = 00010
       -- reg 13
       X"00003402",
       
        -- FIRST SET
        
        
       -- opcode = 00000000000000000, dr = 01110, sa = 00000,  sb = 00001
       -- reg 14
       X"00003801",
       
       -- opcode = 00000000000000000, dr = 01111, sa = 00000,  sb = 00000
       -- reg 15
       X"00003C00",
       
       -- opcode = 00000000000000000, dr = 10000, sa = 00000,  sb = 00011
       -- reg 16
       X"00004003",
       
       -- opcode = 00000000000000000, dr = 10001, sa = 00000,  sb = 00011
       -- reg 17
       X"00004402",
       
       -- opcode = 00000000000000000, dr = 10010, sa = 00000,  sb = 00001
       -- reg 18
       X"00004801",
       
       -- opcode = 00000000000000000, dr = 10011, sa = 00000,  sb = 00000
       -- reg 19
       X"00004C00",
       
       -- opcode = 00000000000000000, dr = 10100, sa = 00000,  sb = 00011
       -- reg 20
       X"00005003",
       
       -- opcode = 00000000000000000, dr = 10101, sa = 00000,  sb = 00010
       -- reg 21
       X"00005402",
       
       -- opcode = 00000000000000000, dr = 10110, sa = 00000,  sb = 00001
       -- reg 22
       X"00005801",
       
       -- opcode = 00000000000000000, dr = 10111, sa = 00000,  sb = 00000
       -- reg 23
       X"00005C00",
       
       -- opcode = 00000000000000000, dr = 11000, sa = 00000,  sb = 00011
       -- reg 24
       X"00006003",
       
       -- opcode = 00000000000000000, dr = 11001, sa = 00000,  sb = 00011
       -- reg 25
       X"00006402",
       
       -- opcode = 00000000000000000, dr = 11010, sa = 00000,  sb = 00001
       -- reg 26
       X"00006801",
       
       -- opcode = 00000000000000000, dr = 11011, sa = 00000,  sb = 00000
       -- reg 27
       X"00006C00",
       
       -- opcode = 00000000000000000, dr = 11100, sa = 00000,  sb = 00011
       -- reg 28
       X"00007003",
       
       -- opcode = 00000000000000000, dr = 11101, sa = 00000,  sb = 00010
       -- reg 29
       X"00007402",
       
       -- opcode = 00000000000000000, dr = 11110, sa = 00000,  sb = 00001
       -- reg 30
       X"00007801",
       
       -- SECOND SET
       
       -- opcode = 00000000000000001, dr = 11111, sa = 00000,  sb = 00000
       -- reg 31
       X"0000FC00",
       
       -- opcode = 00000000000000000, dr = 00000, sa = 00000,  sb = 00011
       -- reg 32
       X"00000003",

       
       -- ADI - Adds reg1 with constant 3 into reg 0
       
       -- opcode = 0000000000000001|0, dr = 000|00, sa = 00|001,  sb = 0|0011
       X"00010023",
       
       
       -- LD - loads value from location 0 (ie the number 0) into reg 2
       
       -- opcode = 0000000000000001|1, dr = 000|10, sa = 00|000,  sb = 0|0000
       X"00018800",
       
       
       -- SR - shift value from reg 3 into reg 4
       
       -- opcode = 0000000000000010|0, dr = 001|00, sa = 00|000,  sb = 0|0011
       X"00021003", 
       
       
       -- INC - increment the value from reg 5 and store in reg 6
       
       -- opcode = 0000000000000010|1, dr = 001|10, sa = 00|101,  sb = 0|0000
       X"000298A0", 
       
       
       -- NOT - not(reg7) and store in reg 8
       
       -- opcode = 0000000000000011|0, dr = 010|00, sa = 00|111,  sb = 0|0000
       X"000320E0",
       
       
       -- ADD - reg 9 + reg 10 into reg 11
       
       -- opcode = 0000000000000011|1, dr = 010|11, sa = 01|001,  sb = 0|1010
       X"0003AD2A",
       
       
       -- unconditional branch
       
       -- opcode = 0000000000000000|0, dr = 000|00, sa = 00|000,  sb = 0|0000
       X"00000000", 
       
       
       -- conditional branch - if not zero reg 12 + reg 13 into reg 14
       
       -- opcode = 0000000000001000|0, dr = 011|10, sa = 01|100,  sb = 0|1101
       X"0008398D", 
       
       
       X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- THIRD SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- FOURTH SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- FIFTH SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- SIXTH SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- SEVENTH SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- EIGHTH SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- NINTH SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- TENTH SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- ELEVENTH SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- TWELFTH SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- THIRTEENTH SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- FOURTEENTH SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- FIFTEENTH SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- SIXTEENTH SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- SEVENTEENTH SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- EIGHTEENTH SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- NINETEENTH SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- TWENTIETH SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- TWENTY FIRST SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- TWENTY SECOND SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- TWENTY THIRD SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- TWENTY FOURTH SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- TWENTY FIFTH SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- TWENTY SIXTH SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- TWENTY SEVENTH SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- TWENTY EIGHTH SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- TWENTY NINTH SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- THIRTIETH SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       
       -- THIRTY FIRST SET
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000",
       X"00000000", X"00000000", X"00000000",X"00000000");
       
    variable addr:integer range 0 to 511;
begin -- the following type conversion function is in std_logic_arith

    addr:= conv_integer(unsigned(address(8 downto 0)));
    
    
    if MW ='1' and clk = '1' then
        data_mem(addr):= write_data;
    elsif MW ='0' and clk ='1' then
        read_data <= data_mem(addr) after 10 ns;
    end if;
    
end process;

end Behavioral;
