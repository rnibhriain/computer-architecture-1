----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 22.12.2020 21:07:02
-- Design Name: 
-- Module Name: control_memory - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity control_memory is
Port (  FL : out std_logic; -- 0
        RZ : out std_logic; -- 1
        RN : out std_logic; -- 2
        RC : out std_logic; -- 3
        RV : out std_logic; -- 4
        
        
        MW : out std_logic; -- 5
        MM : out std_logic; -- 6
        RW : out std_logic; -- 7
        MD : out std_logic; -- 8
        FS : out std_logic_vector(4 downto 0); -- 9 to 13
        MB : out std_logic; -- 14
        
        
        TB : out std_logic; -- 15
        TA : out std_logic; -- 16
        TD : out std_logic; -- 17
        PL : out std_logic; -- 18
        PI : out std_logic; -- 19
        IL : out std_logic; -- 20
        MC : out std_logic; -- 21
        MS : out std_logic_vector(2 downto 0); -- 22 to 24
        NA : out std_logic_vector(16 downto 0); -- 25 to 41
        IN_CAR : in std_logic_vector(16 downto 0));
end control_memory;

architecture Behavioral of control_memory is

    type mem_array is array(0 to 255) of std_logic_vector(41 downto 0);

begin

memory_m: process(IN_CAR)
    variable control_mem : mem_array:= (
    
        -- |41 25|2422|21|20|19|18|17|16|15|14|13 9|8|7|6|5|4|3|2|1|0|
        -- | Next Address | MS | M| I| P| P| T| T| T| M| FS |M|R|M|M|R|R|R|R|F|
        -- | Next Address | MS | C| L| I| L| D| A| B| B| FS |D|W|M|W|V|C|N|Z|L|
        
        -- |41 25|2422|21|20|19|18|17|16|15|14|13 9|8|7|6|5|4|3|2|1|0|
        -- | Next Address    | MS | M| I| P| P| T| T| T| M| FS  |M|R|M|M|R|R|R|R|F|
        -- | Next Address    | MS | C| L| I| L| D| A| B| B| FS  |D|W|M|W|V|C|N|Z|L|
        -- 00000000000000000  001   1  1  1  0  0  0  0  1 00000 0 1 1 0 1 1 1 1 1   
        
        -- reset everything and load values into registers from 0 to 31
        "000000000000000000011110000100000011011111",-- 00
               
        
        -- |41 25|2422|21|20|19|18|17|16|15|14|13 9|8|7|6|5|4|3|2|1|0|
        -- | Next Address    | MS | M| I| P| P| T| T| T| M| FS  |M|R|M|M|R|R|R|R|F|
        -- | Next Address    | MS | C| L| I| L| D| A| B| B| FS  |D|W|M|W|V|C|N|Z|L|
        -- 00000000000000010  001   0  1  1  0  1  1  0  1 00000 0 1 1 0 1 1 1 1 1  
        
        -- load register 32
        "000000000000000100010110110100000011011111",-- 01
        
        -- |41 25|2422|21|20|19|18|17|16|15|14|13 9|8|7|6|5|4|3|2|1|0|
        -- | Next Address    | MS | M| I| P| P| T| T| T| M| FS  |M|R|M|M|R|R|R|R|F|
        -- | Next Address    | MS | C| L| I| L| D| A| B| B| FS  |D|W|M|W|V|C|N|Z|L|
        -- 00000000000000011  000   0  1  1  0  0  0  0  1 00010 0 1 1 0 0 0 0 0 1 
        
        -- ADI
        "000000000000000110000110000100010011000001",-- 02
        
        -- |41 25|2422|21|20|19|18|17|16|15|14|13 9|8|7|6|5|4|3|2|1|0|
        -- | Next Address    | MS | M| I| P| P| T| T| T| M| FS  |M|R|M|M|R|R|R|R|F|
        -- | Next Address    | MS | C| L| I| L| D| A| B| B| FS  |D|W|M|W|V|C|N|Z|L|
        -- 00000000000000100  000   0  1  1  0  0  0  0  0 00000 1 1 1 0 0 0 0 0 1
        
        -- LD
        "000000000000001000000110000000000111000001",-- 03
        
        -- |41 25|2422|21|20|19|18|17|16|15|14|13 9|8|7|6|5|4|3|2|1|0|
        -- | Next Address    | MS | M| I| P| P| T| T| T| M| FS  |M|R|M|M|R|R|R|R|F|
        -- | Next Address    | MS | C| L| I| L| D| A| B| B| FS  |D|W|M|W|V|C|N|Z|L|
        -- 00000000000000100  000   0  1  1  0  0  0  0  1 10100 0 1 1 0 0 0 0 0 1
        
        -- SR
        "000000000000001000000110000110100011000001",-- 04
        
        -- |41 25|2422|21|20|19|18|17|16|15|14|13 9|8|7|6|5|4|3|2|1|0|
        -- | Next Address    | MS | M| I| P| P| T| T| T| M| FS  |M|R|M|M|R|R|R|R|F|
        -- | Next Address    | MS | C| L| I| L| D| A| B| B| FS  |D|W|M|W|V|C|N|Z|L|
        -- 00000000000000101  000   0  1  1  0  0  0  0  1 00001 0 1 1 0 0 0 0 0 1
        
        -- INC 
        "000000000000001010000110000100001011000001",-- 05
        
        -- |41 25|2422|21|20|19|18|17|16|15|14|13 9|8|7|6|5|4|3|2|1|0|
        -- | Next Address    | MS | M| I| P| P| T| T| T| M| FS  |M|R|M|M|R|R|R|R|F|
        -- | Next Address    | MS | C| L| I| L| D| A| B| B| FS  |D|W|M|W|V|C|N|Z|L|
        -- 00000000000000110  000   0  1  1  0  0  0  0  1 01110 0 1 1 0 0 0 0 0 1
        
        -- NOT
        "000000000000001100000110000101110011000001",-- 06
        
        -- |41 25|2422|21|20|19|18|17|16|15|14|13 9|8|7|6|5|4|3|2|1|0|
        -- | Next Address    | MS | M| I| P| P| T| T| T| M| FS  |M|R|M|M|R|R|R|R|F|
        -- | Next Address    | MS | C| L| I| L| D| A| B| B| FS  |D|W|M|W|V|C|N|Z|L|
        -- 00000000000000111  000   0  1  1  0  0  0  0  0 00010 0 1 1 0 0 0 0 0 1
        
        -- ADD
        "000000000000000000000000000000000000000000",-- 07
        
        -- |41 25|2422|21|20|19|18|17|16|15|14|13 9|8|7|6|5|4|3|2|1|0|
        -- | Next Address    | MS | M| I| P| P| T| T| T| M| FS  |M|R|M|M|R|R|R|R|F|
        -- | Next Address    | MS | C| L| I| L| D| A| B| B| FS  |D|W|M|W|V|C|N|Z|L|
        -- 00000000000010000  001   0  1  1  0  0  0  0  0 00000 0 0 1 0 0 0 0 0 0
        
        -- unconditional jump
        "000000000000100000010110000000000001000000",-- 08
        
        
        
        
        "000000000000000000000000000000000000000000",-- 09
        "000000000000000000000000000000000000000000",-- 0A
        "000000000000000000000000000000000000000000",-- 0B
        "000000000000000000000000000000000000000000",-- 0C
        "000000000000000000000000000000000000000000",-- 0D
        "000000000000000000000000000000000000000000",-- 0E
        "000000000000000000000000000000000000000000",-- 0F
        
        
        -- |41 25|2422|21|20|19|18|17|16|15|14|13 9|8|7|6|5|4|3|2|1|0|
        -- | Next Address    | MS | M| I| P| P| T| T| T| M| FS  |M|R|M|M|R|R|R|R|F|
        -- | Next Address    | MS | C| L| I| L| D| A| B| B| FS  |D|W|M|W|V|C|N|Z|L|
        -- 00000000011000000  111   0  1  1  0  0  0  0  0 00010 0 0 1 0 0 0 0 0 1
        
        -- conditional branch if not zero
        "000000000110000001110110000000010001000001",-- 10
        
        
        
        "000000000000000000000000000000000000000000",-- 11
        "000000000000000000000000000000000000000000",-- 12
        "000000000000000000000000000000000000000000",-- 13
        "000000000000000000000000000000000000000000",-- 14
        "000000000000000000000000000000000000000000",-- 15
        "000000000000000000000000000000000000000000",-- 16
        "000000000000000000000000000000000000000000",-- 17
        
        "000000000000000000000000000000000000000000",-- 18
        "000000000000000000000000000000000000000000",-- 19
        "000000000000000000000000000000000000000000",-- 1A
        "000000000000000000000000000000000000000000",-- 1B
        "000000000000000000000000000000000000000000",-- 1C
        "000000000000000000000000000000000000000000",-- 1D
        "000000000000000000000000000000000000000000",-- 1E
        "000000000000000000000000000000000000000000",-- 1F
        
        "000000000000000000000000000000000000000000",-- 20
        "000000000000000000000000000000000000000000",-- 21
        "000000000000000000000000000000000000000000",-- 22
        "000000000000000000000000000000000000000000",-- 23
        "000000000000000000000000000000000000000000",-- 24
        "000000000000000000000000000000000000000000",-- 25
        "000000000000000000000000000000000000000000",-- 26
        "000000000000000000000000000000000000000000",-- 27
        
        "000000000000000000000000000000000000000000",-- 28
        "000000000000000000000000000000000000000000",-- 29
        "000000000000000000000000000000000000000000",-- 2A
        "000000000000000000000000000000000000000000",-- 2B
        "000000000000000000000000000000000000000000",-- 2C
        "000000000000000000000000000000000000000000",-- 2D
        "000000000000000000000000000000000000000000",-- 2E
        "000000000000000000000000000000000000000000",-- 2F
        
        
        "000000000000000000000000000000000000000000",-- 30
        "000000000000000000000000000000000000000000",-- 31
        "000000000000000000000000000000000000000000",-- 32
        "000000000000000000000000000000000000000000",-- 33
        "000000000000000000000000000000000000000000",-- 34
        "000000000000000000000000000000000000000000",-- 35
        "000000000000000000000000000000000000000000",-- 36
        "000000000000000000000000000000000000000000",-- 37
        
        "000000000000000000000000000000000000000000",-- 38
        "000000000000000000000000000000000000000000",-- 39
        "000000000000000000000000000000000000000000",-- 3A
        "000000000000000000000000000000000000000000",-- 3B
        "000000000000000000000000000000000000000000",-- 3C
        "000000000000000000000000000000000000000000",-- 3D
        "000000000000000000000000000000000000000000",-- 3E
        "000000000000000000000000000000000000000000",-- 3F
        
        
        "000000000000000000000000000000000000000000",-- 40
        "000000000000000000000000000000000000000000",-- 41
        "000000000000000000000000000000000000000000",-- 42
        "000000000000000000000000000000000000000000",-- 43
        "000000000000000000000000000000000000000000",-- 44
        "000000000000000000000000000000000000000000",-- 45
        "000000000000000000000000000000000000000000",-- 46
        "000000000000000000000000000000000000000000",-- 47
        
        "000000000000000000000000000000000000000000",-- 48
        "000000000000000000000000000000000000000000",-- 49
        "000000000000000000000000000000000000000000",-- 4A
        "000000000000000000000000000000000000000000",-- 4B
        "000000000000000000000000000000000000000000",-- 4C
        "000000000000000000000000000000000000000000",-- 4D
        "000000000000000000000000000000000000000000",-- 4E
        "000000000000000000000000000000000000000000",-- 4F
        
        
        
        "000000000000000000000000000000000000000000",-- 50
        "000000000000000000000000000000000000000000",-- 51
        "000000000000000000000000000000000000000000",-- 52
        "000000000000000000000000000000000000000000",-- 53
        "000000000000000000000000000000000000000000",-- 54
        "000000000000000000000000000000000000000000",-- 55
        "000000000000000000000000000000000000000000",-- 56
        "000000000000000000000000000000000000000000",-- 57
        
        "000000000000000000000000000000000000000000",-- 58
        "000000000000000000000000000000000000000000",-- 59
        "000000000000000000000000000000000000000000",-- 5A
        "000000000000000000000000000000000000000000",-- 5B
        "000000000000000000000000000000000000000000",-- 5C
        "000000000000000000000000000000000000000000",-- 5D
        "000000000000000000000000000000000000000000",-- 5E
        "000000000000000000000000000000000000000000",-- 5F
        
        
        
        "000000000000000000000000000000000000000000",-- 60
        "000000000000000000000000000000000000000000",-- 61
        "000000000000000000000000000000000000000000",-- 62
        "000000000000000000000000000000000000000000",-- 63
        "000000000000000000000000000000000000000000",-- 64
        "000000000000000000000000000000000000000000",-- 65
        "000000000000000000000000000000000000000000",-- 66
        "000000000000000000000000000000000000000000",-- 67
        
        "000000000000000000000000000000000000000000",-- 68
        "000000000000000000000000000000000000000000",-- 69
        "000000000000000000000000000000000000000000",-- 6A
        "000000000000000000000000000000000000000000",-- 6B
        "000000000000000000000000000000000000000000",-- 6C
        "000000000000000000000000000000000000000000",-- 6D
        "000000000000000000000000000000000000000000",-- 6E
        "000000000000000000000000000000000000000000",-- 6F
        
        
        
        "000000000000000000000000000000000000000000",-- 70
        "000000000000000000000000000000000000000000",-- 71
        "000000000000000000000000000000000000000000",-- 72
        "000000000000000000000000000000000000000000",-- 73
        "000000000000000000000000000000000000000000",-- 74
        "000000000000000000000000000000000000000000",-- 75
        "000000000000000000000000000000000000000000",-- 76
        "000000000000000000000000000000000000000000",-- 77
        
        "000000000000000000000000000000000000000000",-- 78
        "000000000000000000000000000000000000000000",-- 79
        "000000000000000000000000000000000000000000",-- 7A
        "000000000000000000000000000000000000000000",-- 7B
        "000000000000000000000000000000000000000000",-- 7C
        "000000000000000000000000000000000000000000",-- 7D
        "000000000000000000000000000000000000000000",-- 7E
        "000000000000000000000000000000000000000000",-- 7F
        
        
        "000000000000000000000000000000000000000000",-- 80
        "000000000000000000000000000000000000000000",-- 81
        "000000000000000000000000000000000000000000",-- 82
        "000000000000000000000000000000000000000000",-- 83
        "000000000000000000000000000000000000000000",-- 84
        "000000000000000000000000000000000000000000",-- 85
        "000000000000000000000000000000000000000000",-- 86
        "000000000000000000000000000000000000000000",-- 87
        
        "000000000000000000000000000000000000000000",-- 88
        "000000000000000000000000000000000000000000",-- 89
        "000000000000000000000000000000000000000000",-- 8A
        "000000000000000000000000000000000000000000",-- 8B
        "000000000000000000000000000000000000000000",-- 8C
        "000000000000000000000000000000000000000000",-- 8D
        "000000000000000000000000000000000000000000",-- 8E
        "000000000000000000000000000000000000000000",-- 8F
        
        
        
        "000000000000000000000000000000000000000000",-- 90
        "000000000000000000000000000000000000000000",-- 91
        "000000000000000000000000000000000000000000",-- 92
        "000000000000000000000000000000000000000000",-- 93
        "000000000000000000000000000000000000000000",-- 94
        "000000000000000000000000000000000000000000",-- 95
        "000000000000000000000000000000000000000000",-- 96
        "000000000000000000000000000000000000000000",-- 97
        
        "000000000000000000000000000000000000000000",-- 98
        "000000000000000000000000000000000000000000",-- 99
        "000000000000000000000000000000000000000000",-- 9A
        "000000000000000000000000000000000000000000",-- 9B
        "000000000000000000000000000000000000000000",-- 9C
        "000000000000000000000000000000000000000000",-- 9D
        "000000000000000000000000000000000000000000",-- 9E
        "000000000000000000000000000000000000000000",-- 9F
        
        
        
        "000000000000000000000000000000000000000000",-- A0
        "000000000000000000000000000000000000000000",-- A1
        "000000000000000000000000000000000000000000",-- A2
        "000000000000000000000000000000000000000000",-- A3
        "000000000000000000000000000000000000000000",-- A4
        "000000000000000000000000000000000000000000",-- A5
        "000000000000000000000000000000000000000000",-- A6
        "000000000000000000000000000000000000000000",-- A7
        
        "000000000000000000000000000000000000000000",-- A8
        "000000000000000000000000000000000000000000",-- A9
        "000000000000000000000000000000000000000000",-- AA
        "000000000000000000000000000000000000000000",-- AB
        "000000000000000000000000000000000000000000",-- AC
        "000000000000000000000000000000000000000000",-- AD
        "000000000000000000000000000000000000000000",-- AE
        "000000000000000000000000000000000000000000",-- AF
        
        
        
        "000000000000000000000000000000000000000000",-- B0
        "000000000000000000000000000000000000000000",-- B1
        "000000000000000000000000000000000000000000",-- B2
        "000000000000000000000000000000000000000000",-- B3
        "000000000000000000000000000000000000000000",-- B4
        "000000000000000000000000000000000000000000",-- B5
        "000000000000000000000000000000000000000000",-- B6
        "000000000000000000000000000000000000000000",-- B7
        
        "000000000000000000000000000000000000000000",-- B8
        "000000000000000000000000000000000000000000",-- B9
        "000000000000000000000000000000000000000000",-- BA
        "000000000000000000000000000000000000000000",-- BB
        "000000000000000000000000000000000000000000",-- BC
        "000000000000000000000000000000000000000000",-- BD
        "000000000000000000000000000000000000000000",-- BE
        "000000000000000000000000000000000000000000",-- BF
        
        -- |41 25|2422|21|20|19|18|17|16|15|14|13 9|8|7|6|5|4|3|2|1|0|
        -- | Next Address    | MS | M| I| P| P| T| T| T| M| FS  |M|R|M|M|R|R|R|R|F|
        -- | Next Address    | MS | C| L| I| L| D| A| B| B| FS  |D|W|M|W|V|C|N|Z|L|
        -- 00000000011000001  000   0  1  0  0  0  0  0  0 00000 0 0 1 0 0 0 0 0 0
        
        -- If Fetching
        "000000000110000010000100000000000001000000",-- C0
        
        -- |41 25|2422|21|20|19|18|17|16|15|14|13 9|8|7|6|5|4|3|2|1|0|
        -- | Next Address    | MS | M| I| P| P| T| T| T| M| FS  |M|R|M|M|R|R|R|R|F|
        -- | Next Address    | MS | C| L| I| L| D| A| B| B| FS  |D|W|M|W|V|C|N|Z|L|
        -- 00000000000000000  001   1  0  0  0  0  0  0  0 00000 0 1 0 0 0 0 0 0 0
        
        -- Exiting
        "000000000000000000011000000000000010000000",-- C1
        "000000000000000000000000000000000000000000",-- C2
        "000000000000000000000000000000000000000000",-- C3
        "000000000000000000000000000000000000000000",-- C4
        "000000000000000000000000000000000000000000",-- C5
        "000000000000000000000000000000000000000000",-- C6
        "000000000000000000000000000000000000000000",-- C7
        
        "000000000000000000000000000000000000000000",-- C8
        "000000000000000000000000000000000000000000",-- C9
        "000000000000000000000000000000000000000000",-- CA
        "000000000000000000000000000000000000000000",-- CB
        "000000000000000000000000000000000000000000",-- CC
        "000000000000000000000000000000000000000000",-- CD
        "000000000000000000000000000000000000000000",-- CE
        "000000000000000000000000000000000000000000",-- CF
        
        
        "000000000000000000000000000000000000000000",-- D0
        "000000000000000000000000000000000000000000",-- D1
        "000000000000000000000000000000000000000000",-- D2
        "000000000000000000000000000000000000000000",-- D3
        "000000000000000000000000000000000000000000",-- D4
        "000000000000000000000000000000000000000000",-- D5
        "000000000000000000000000000000000000000000",-- D6
        "000000000000000000000000000000000000000000",-- D7
       
        "000000000000000000000000000000000000000000",-- D8
        "000000000000000000000000000000000000000000",-- D9
        "000000000000000000000000000000000000000000",-- DA
        "000000000000000000000000000000000000000000",-- DB
        "000000000000000000000000000000000000000000",-- DC
        "000000000000000000000000000000000000000000",-- DD
        "000000000000000000000000000000000000000000",-- DE
        "000000000000000000000000000000000000000000",-- DF
        
        
        "000000000000000000000000000000000000000000",-- E0
        "000000000000000000000000000000000000000000",-- E1
        "000000000000000000000000000000000000000000",-- E2
        "000000000000000000000000000000000000000000",-- E3
        "000000000000000000000000000000000000000000",-- E4
        "000000000000000000000000000000000000000000",-- E5
        "000000000000000000000000000000000000000000",-- E6
        "000000000000000000000000000000000000000000",-- E7
        
        "000000000000000000000000000000000000000000",-- E8
        "000000000000000000000000000000000000000000",-- E9
        "000000000000000000000000000000000000000000",-- EA
        "000000000000000000000000000000000000000000",-- EB
        "000000000000000000000000000000000000000000",-- EC
        "000000000000000000000000000000000000000000",-- ED
        "000000000000000000000000000000000000000000",-- EE
        "000000000000000000000000000000000000000000",-- EF
        
        
        "000000000000000000000000000000000000000000",-- F0
        "000000000000000000000000000000000000000000",-- F1
        "000000000000000000000000000000000000000000",-- F2
        "000000000000000000000000000000000000000000",-- F3
        "000000000000000000000000000000000000000000",-- F4
        "000000000000000000000000000000000000000000",-- F5
        "000000000000000000000000000000000000000000",-- F6
        "000000000000000000000000000000000000000000",-- F7
        
        "000000000000000000000000000000000000000000",-- F8
        "000000000000000000000000000000000000000000",-- F9
        "000000000000000000000000000000000000000000",-- FA
        "000000000000000000000000000000000000000000",-- FB
        "000000000000000000000000000000000000000000",-- FC
        "000000000000000000000000000000000000000000",-- FD
        "000000000000000000000000000000000000000000",-- FE
        "000000000000000000000000000000000000000000" -- FF
    );
    
variable addr : integer range 0 to 255;
variable control_out : std_logic_vector(41 downto 0);

begin
    addr := conv_integer(unsigned(IN_CAR(7 downto 0)));
    control_out := control_mem(addr);
    FL <= control_out(0);
    RZ <= control_out(1);
    RN <= control_out(2);
    RC <= control_out(3);
    RV <= control_out(4);
    
    MW <= control_out(5);
    MM <= control_out(6);
    RW <= control_out(7);
    MD <= control_out(8);
    FS <= control_out(13 downto 9);
    MB <= control_out(14);
    
    TB <= control_out(15);
    TA <= control_out(16);
    TD <= control_out(12);
    PL <= control_out(17);
    PI <= control_out(19);
    IL <= control_out(20);
    MC <= control_out(21);
    MS <= control_out(24 downto 22);
    NA <= control_out(41 downto 25);
    
end process;

end Behavioral;
